
/*
	Is a combinational circuit
	Decides for each pixel what color should be on the screen
	
	Glyph graphics - break the screen into chunks
*/
module BitGen (
	input bright,
	input [7:0] pixelData,
	input [9:0] hCount, vCount,
	output reg [7:0] rgb);
	

endmodule
