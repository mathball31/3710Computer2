
module BitGen ();

endmodule
