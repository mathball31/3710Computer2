
module VGAcontrol ();

/* 50MHz clock with 60 fps (60Hz frame rate) */

endmodule
